Switch testbench

.param L = 0.18U
.param WL = 3
.param W = { WL * L}

.param Vdd = 1.8
.param Vg = Vdd

VDD 1 0 dc Vdd
VGG 2 0 dc Vg

MN1 1 2 0 0 NMOS L=L W=W

.dc VGG 0 Vg 0.01

.plot gm(MN1)

.include p18_model_card.inc
.include p18_cmos_models_ss.inc