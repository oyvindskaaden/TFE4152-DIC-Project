//
//
// Top-level verilog module example
//

module re_control(Expose, Erase, ADC, NRE_1, NRE_2,
	Init, Exp_increase, Exp_decrease, Reset, Clk);

	input Init, Exp_increase, Exp_decrease, Reset, Clk;
	output Expose, Erase, ADC, NRE_1, NRE_2;
	
	
	//
	// Your code goes here
	//
	
endmodule // re_control

