module FSM_ex_control(
	input 	logic 			clk;
	input 	logic 			reset;
	input 	logic 			init;
	input 	wire 				ex_done;
	output 	wire 				ex_start;

	output 	wire [1:0] 	nre;
	output 	wire 				adc;
	output 	wire 				expose;
	output 	wire 				erase;
);



endmodule