module FSM_ex_control(
	input logic clk;
	input logic reset;
	input logic init;
	output wire ex_start;
	input wire ex_done;
);



endmodule